module aa;
wire signed [4:-4] a;
assign a=2%4;
endmodule 
